  // ls
 repeat (10)
abc;
