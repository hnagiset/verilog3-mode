   /*
The quick brown fox
  module
*/
  // basic-test.sv
// hello
   module hello();
abc;
def;
   module hello();
abc;
     if (abc)
       if (abc)
def;
       else
         begin
         ghi;
         ghi;
  `ifdef hi
           if abc
             `endif
             afunction(a,
                   b,
                   c);
             bfunction(
a,
             cfunction(
  a,
  a,
  a,
  a)
                   b, c);
           while (a)
xyz;
         ghi;
         ghi;
           end
while (a) begin
 abc;
end

     fork;
       ab;
     join

     wait fork;
      ab;
xyz;
def;
   module hello();
abc;
def;
endmodule
endmodule
endmodule
