module hello();
abc;
def;
endmodule
