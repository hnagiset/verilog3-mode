
function hi();
function hi();
abc;
  extern function hi();
  externa function hi();
    a;
    endfunction
  import function hi();
  pure virtual function hi();
  virtual function hi();
abc;
endfunction
abc;
endfunction
endfunction
